--
-- VHDL Architecture Temperature_PIDcontroller_lib.tempeerature_model.Behavioral
--
-- Created:
--          by - Abdelaziz.UNKNOWN (ABDULLAH)
--          at - 14:40:01 05/ 1/2025
--
-- using Mentor Graphics HDL Designer(TM) 2018.2 (Build 19)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY temperature_model IS
  port (
        clk             : in  std_logic;
        reset           : in  std_logic;
        fan_speed_in    : in  integer range 0 to 100;
        ambient_temp_in : in  integer range 0 to 100;  -- Ambient temperature
        current_temp_out: out integer range 0 to 100
    );
END ENTITY temperature_model;

--
ARCHITECTURE Behavioral OF temperature_model IS
  
   -- Internal signals
    signal internal_temp      : real := 25.0;  -- Using 'real' for better precision
    signal prev_temp          : real := 25.0;
    signal delta_temp         : real := 0.0;
    signal normalized_fan_speed: real := 0.0;

    -- Constants
    constant thermal_resistance : real := 2.0;  -- Adjust as needed (how much temp rises per unit heat)
    constant thermal_capacitance: real := 0.1;  -- Adjust (how much the FPGA resists temp change)
    constant fpga_heat_generation : real := 1.0; -- Base heat generated by FPGA 


BEGIN
  process (clk, reset)
    begin
        if reset = '0' then
            internal_temp <= 25.0;
            prev_temp <= 25.0;
            current_temp_out <= 25;
        elsif rising_edge(clk) then

            -- Normalize fan speed and make it non-linear
            normalized_fan_speed <= real(fan_speed_in) / 100.0;
            normalized_fan_speed <= normalized_fan_speed * normalized_fan_speed; -- Non-linear curve

            -- Calculate temperature change (simplified heat transfer)
            delta_temp <= (fpga_heat_generation - (internal_temp - real(ambient_temp_in)) / thermal_resistance - normalized_fan_speed * (internal_temp - real(ambient_temp_in)) / thermal_resistance) * thermal_capacitance;

            -- Apply thermal inertia (temperature doesn't change instantly)
            internal_temp <= internal_temp + delta_temp;

            -- Keep temperature within bounds
            if internal_temp > 100.0 then
                internal_temp <= 100.0;
            elsif internal_temp < 0.0 then
                internal_temp <= 0.0;
            end if;

            current_temp_out <= integer(internal_temp); -- Output as integer

            prev_temp <= internal_temp;

        end if;
    end process;
END ARCHITECTURE Behavioral;

